module  PipelineCPU (resetn,clock,
					operand0, operand1,
					hex0, hex1, hex2, hex3, hex4, hex5, hex6, hex7, led0, led1, led);
//���嶥��ģ�� pipelined_computer����Ϊ�����ļ��Ķ�����ڣ���ͼ 1-1 ��������ʱָ���� 

	input [7:0] operand0;
	input [3:0]  operand1;
	//input [3:0] operand0, operand1;
	output [6:0] hex0, hex1, hex2, hex3, hex4, hex5, hex6, hex7;
	output [3:0] led0, led1;
	output led;
	wire [31:0] in_port0,in_port1,out_port0,out_port1;
	wire [6:0] hex_null;
	wire mem_dataout, io_read_data;
	
	assign in_port0 = {24'b0, operand0[7:0]};
	assign in_port1 = {24'b0, 8'b11001010};
	//operand_to_in_port binary32_operand0(mem_clock, operand0, in_port0);
    //operand_to_in_port binary32_operand1(mem_clock, operand1, in_port1);
    
    //binary_to_sevenseg LED8_in_port0(mem_clock, in_port0, hex7, hex6);
    //binary_to_sevenseg LED8_in_port1(mem_clock, in_port1, hex5, hex4);
	
    binary_to_sevenseg LED8_out_port0(mem_clock, out_port0, hex_null, hex3);
    
    assign hex0 = 7'b111_1111;
    assign hex1 = 7'b111_1111;
    assign hex2 = 7'b111_1111;
    assign hex4 = 7'b111_1111;
    assign hex5 = 7'b111_1111;
    assign hex6 = 7'b111_1111;
    assign hex7 = 7'b111_1111;
    //assign led0 = operand0;
    //assign led1 = operand1;
    assign led = ~resetn;
    //insert I/O
	
	input          resetn, clock; 
//������������� module ����罻���������źţ�������λ�ź� resetn��ʱ���ź� clock�� 
//�Լ�һ���� clock ͬƵ�ʵ������ mem_clock �źš�mem_clock ����ָ��ͬ�� ROM �� 
//����ͬ�� RAM ʹ�ã��䲨����Ҫ�б���ʵ��һ�� 
//��Щ�źſ�������������֤ʱ������۲��źš� 
	wire  [31:0]  pc,ealu,malu,walu; 
	//output  [31:0]  pc,inst,ealu,malu,walu,da,db, wpcir; 
//ģ�����ڷ�������Ĺ۲��źš�ȱʡΪ wire �͡� 
	wire   [31:0]  bpc,jpc,npc,pc4,ins, inst;     
//ģ��以���������ݻ������Ϣ���ź���,��Ϊ 32 λ���źš�IF ȡָ��׶Ρ� 
	wire   [31:0]  dpc4,da,db,dimm; 
//ģ��以���������ݻ������Ϣ���ź���,��Ϊ 32 λ���źš�ID ָ������׶Ρ� 
	wire   [31:0]  epc4,ea,eb,eimm;  
//ģ��以���������ݻ������Ϣ���ź���,��Ϊ 32 λ���źš�EXE ָ������׶Ρ� 
	wire   [31:0]  mb,mmo; 
//ģ��以���������ݻ������Ϣ���ź���,��Ϊ 32 λ���źš�MEM �������ݽ׶Ρ� 
	wire   [31:0]  wmo,wdi; 
//ģ��以���������ݻ������Ϣ���ź���,��Ϊ 32 λ���źš�WB ��д�Ĵ����׶Ρ� 
	wire   [4:0]   drn,ern0,ern,mrn,wrn; 
//ģ��以����ͨ����ˮ�߼Ĵ������ݽ���Ĵ����ŵ��ź��ߣ��Ĵ����ţ�32 ����Ϊ 5bit�� 
	wire   [3:0]   daluc,ealuc; 
//ID �׶��� EXE �׶�ͨ����ˮ�߼Ĵ������ݵ� aluc �����źţ�4bit�� 
	wire   [1:0]   pcsource; 
//CU ģ���� IF �׶�ģ�鴫�ݵ� PC ѡ���źţ�2bit�� 
	wire          wpcir; 
// CU ģ�鷢���Ŀ�����ˮ��ͣ�ٵĿ����źţ�ʹ PC �� IF/ID ��ˮ�߼Ĵ������ֲ��䡣 
	wire          dwreg,dm2reg,dwmem,daluimm,dshift,djal;  // id stage 
// ID �׶β���������������ˮ���������źš� 
	wire          ewreg,em2reg,ewmem,ealuimm,eshift,ejal;  // exe stage 
//������ ID/EXE ��ˮ�߼Ĵ�����EXE �׶�ʹ�ã�����Ҫ��������ˮ���������źš� 
	wire          mwreg,mm2reg,mwmem;  // mem stage 
//������ EXE/MEM ��ˮ�߼Ĵ�����MEM �׶�ʹ�ã�����Ҫ��������ˮ���������źš�       
	wire          wwreg,wm2reg;          // wb stage 
//������ MEM/WB ��ˮ�߼Ĵ�����WB �׶�ʹ�õ��źš� 
	
	wire mem_clock;
	assign mem_clock = ~clock;
	
	pipepc  prog_cnt ( npc,wpcir,clock,resetn,pc ); //���������ģ�飬����ǰ��һ�� IF ��ˮ�ε����롣       
	pipeif  if_stage   ( pcsource,pc,bpc,da,jpc,npc,pc4,ins,mem_clock );  //  IF stage 
//IF ȡָ��ģ�飬ע�����а�����ָ��ͬ�� ROM �洢����ͬ���źţ� 
//���������ģ��� mem_clock �źţ�ģ���ڶ���Ϊ rom_clk��
//ע�� mem_clock�� 
//ʵ���пɲ���ϵͳ clock �ķ����ź���Ϊ mem_clock���༴ rom_clock��, 
//�������źŰ�����ĵĴ���ʱ�䡣 
	pipeir  inst_reg   ( pc4,ins,wpcir,clock,resetn,dpc4,inst );        // IF/ID ��ˮ�߼Ĵ��� 
//IF/ID ��ˮ�߼Ĵ���ģ�飬��н� IF �׶κ� ID �׶ε���ˮ���� 
//�� clock ������ʱ���� IF �׶��贫�ݸ� ID �׶ε���Ϣ�������� IF/ID ��ˮ�߼Ĵ��� 
//�У��������� ID �׶Ρ�       
	pipeid  id_stage  ( mwreg,mrn,ern,ewreg,em2reg,mm2reg,dpc4,inst,
	                    wrn,wdi,ealu,malu,mmo,wwreg,mem_clock,resetn,
	                    bpc,jpc,pcsource,wpcir,dwreg,dm2reg,dwmem,daluc,
	                    daluimm,da,db,dimm,drn,dshift,djal);        //  ID stage 
//ID ָ������ģ�顣ע�����а��������� CU���Ĵ����ѡ��������·���ȡ� 
//���еļĴ����ѣ�����ϵͳ clock �����ؽ��мĴ���д�룬Ҳ���Ǹ��źŴ� WB �׶� 
//����������а�� clock ���ӳ�ʱ�䣬�༴ȷ���ź��ȶ��� 
//�ý׶� CU �����ġ�Ҫ��������ˮ�ߺ󼶵��źŽ϶ࡣ       
	pipedereg  de_reg  ( dwreg,dm2reg,dwmem,daluc,daluimm,da,db,dimm,drn,dshift,
	                     djal,dpc4,clock,resetn,ewreg,em2reg,ewmem,ealuc,ealuimm,
	                     ea,eb,eimm,ern0,eshift,ejal,epc4 );          // ID/EXE ��ˮ�߼Ĵ��� 
//ID/EXE ��ˮ�߼Ĵ���ģ�飬��н� ID �׶κ� EXE �׶ε���ˮ���� 
//�� clock ������ʱ���� ID �׶��贫�ݸ� EXE �׶ε���Ϣ�������� ID/EXE ��ˮ�� 
//�Ĵ����У��������� EXE �׶Ρ�                               
	pipeexe  exe_stage ( ealuc,ealuimm,ea,eb,eimm,eshift,ern0,epc4,ejal,ern,ealu );  // EXE stage        
//EXE ����ģ�顣���а��� ALU �������·���ȡ�                                                 
	pipeemreg  em_reg  ( ewreg,em2reg,ewmem,ealu,eb,ern,clock,resetn,
                         mwreg,mm2reg,mwmem,malu,mb,mrn); // EXE/MEM ��ˮ�߼Ĵ��� 
//EXE/MEM ��ˮ�߼Ĵ���ģ�飬��н� EXE �׶κ� MEM �׶ε���ˮ���� 
//�� clock ������ʱ���� EXE �׶��贫�ݸ� MEM �׶ε���Ϣ�������� EXE/MEM 
//��ˮ�߼Ĵ����У��������� MEM �׶Ρ�      

	pipemem  mem_stage ( mwmem,malu,mb,mem_clock,mmo,
						resetn, out_port0,out_port1,in_port0,in_port1,mem_dataout,io_read_data );        //  MEM stage 
//MEM ���ݴ�ȡģ�顣���а���������ͬ�� RAM �Ķ�д���ʡ�
//ע�� mem_clock�� 
//�������ͬ�� RAM �� mem_clock �źţ�ģ���ڶ���Ϊ ram_clk�� 
//ʵ���пɲ���ϵͳ clock �ķ����ź���Ϊ mem_clock �źţ��༴ ram_clk��, 
//�������źŰ�����ĵĴ���ʱ�䣬Ȼ���� mem_clock ����ʱ�����������д���롣  
    
	pipemwreg  mw_reg  ( mwreg,mm2reg,mmo,malu,mrn,clock,resetn,
                         wwreg,wm2reg,wmo,walu,wrn);     //  MEM/WB ��ˮ�߼Ĵ��� 
//MEM/WB ��ˮ�߼Ĵ���ģ�飬��н� MEM �׶κ� WB �׶ε���ˮ���� 
//�� clock ������ʱ���� MEM �׶��贫�ݸ� WB �׶ε���Ϣ�������� MEM/WB 
//��ˮ�߼Ĵ����У��������� WB �׶Ρ�       
	mux2x32  wb_stage  ( walu,wmo,wm2reg,wdi );          //  WB stage 
//WB д�ؽ׶�ģ�顣��ʵ�ϣ������ԭ��ͼ�Ͽ��Կ������ý׶ε��߼����ܲ���ֻ 
//����һ����·�������Կ��Խ���һ����·����ʵ������ʵ�ָò��֡� 
//��Ȼ�����ר��дһ��������ģ��Ҳ�Ǻܺõġ� 
endmodule

module operand_to_in_port(clk, operand, in_port);
	input clk;
	input [3:0] operand;
	output in_port;
	reg [31:0] in_port;
	
	always @ (posedge clk)
		begin
			in_port <= {28'b0, operand[3:0]};
		end
endmodule

module binary_to_sevenseg(clk, binary, ledsegments0, ledsegments1);
	input clk;
	input [31:0] binary;
	output ledsegments0, ledsegments1;
	reg [6:0] ledsegments0, ledsegments1;
	reg [3:0] Hundreds, Tens, Ones;
	
	integer i;
	always @ (posedge clk)
	begin
		Hundreds = 4'd0;
		Tens = 4'd0;
		Ones = 4'd0;
		
		for (i = 7; i >= 0; i = i - 1)
		begin
			if (Hundreds >= 5)
				Hundreds = Hundreds + 3;
			if (Tens >= 5)
				Tens = Tens + 3;
			if (Ones >= 5)
				Ones = Ones + 3;
				
			Hundreds = Hundreds << 1;
			Hundreds[0] = Tens[3];
			Tens = Tens << 1;
			Tens[0] = Ones[3];
			Ones = Ones << 1;
			Ones[0] = binary[i];
		end
		case (Tens)
			0:ledsegments0 = 7'b100_0000;
			1:ledsegments0 = 7'b111_1001;
			2:ledsegments0 = 7'b010_0100;
			3:ledsegments0 = 7'b011_0000;
			4:ledsegments0 = 7'b001_1001;
			5:ledsegments0 = 7'b001_0010;
			6:ledsegments0 = 7'b000_0010;
			7:ledsegments0 = 7'b111_1000;
			8:ledsegments0 = 7'b000_0000;
			9:ledsegments0 = 7'b001_0000;
			default:ledsegments0 = 7'b111_1111;
		endcase
		case (Ones)
			0:ledsegments1 = 7'b100_0000;
			1:ledsegments1 = 7'b111_1001;
			2:ledsegments1 = 7'b010_0100;
			3:ledsegments1 = 7'b011_0000;
			4:ledsegments1 = 7'b001_1001;
			5:ledsegments1 = 7'b001_0010;
			6:ledsegments1 = 7'b000_0010;
			7:ledsegments1 = 7'b111_1000;
			8:ledsegments1 = 7'b000_0000;
			9:ledsegments1 = 7'b001_0000;
			default:ledsegments1 = 7'b111_1111;
		endcase
	end
endmodule